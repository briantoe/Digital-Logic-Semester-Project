module test_counter:	initial begin			endendmodule