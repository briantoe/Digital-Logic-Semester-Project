module test ();

system #(.debug(1), .program("mem/gcd.mem")) system_test ();

endmodule
