module test ();

system #(.debug(1), .program("mem/example.mem")) system_test ();

endmodule
