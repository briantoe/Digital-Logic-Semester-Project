module counter(out, load, load_data, clk):
	input wire clk;
	output wire[0:15] out;
	input wire load;
	input wire [0:15] load_data;
	
	
	
endmodule