module test ();

system #(.debug(1), .program("src/test/example.mem")) system_test ();

endmodule
