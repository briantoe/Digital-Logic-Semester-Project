module test ();

system #(.debug(1), .file("src/test/example.mem")) system_test ();

endmodule
